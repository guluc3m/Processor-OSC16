--Libraries
library IEEE;
use IEEE.std_logic_1164.all;

--Definition if the entity
entity Processor16Bits is
	port(
		clk: in std_logic;
		rst: in std_logic);
end Processor16Bits;

--Architecture
architecture Behavioral of Processor16Bits is
begin

--cpu : entity work.cpu
	--port map();

--VGA controller
--Keyboard driver
--Main clock process
--Clock divisors processes
end Behavioral;