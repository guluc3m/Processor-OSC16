--Libraries
library IEEE;
use IEEE.std_logic_1164.all;

--Definition if the entity
entity Computer16Bit is
	port(
		clk: in std_logic;
		rst: in std_logic);
end Computer16Bit;

--Architecture
architecture Behavioral of Computer16Bit is
begin

--cpu : entity work.cpu
	--port map();

--VGA controller
--Keyboard driver
--Main clock process
--Clock divisors processes
end Behavioral;